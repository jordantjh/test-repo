module reg_16 (input logic Clk, Reset, Ld_B, Shift_En ,Shift_In, Ld_A,
                      input  logic [7:0]  Ain,Bin, 
                      output logic Shift_Out,
                      output logic [7:0]  Aout,Bout);

		logic A_shift_out;

		reg_8 shift_reg_A (.*, .Shift_In(Shift_In), .Load(Ld_A), .Shift_Out(A_shift_out), .D(Ain), .A(Aout));
		
		reg_8 shift_reg_B (.*, .Reset(0) ,.Shift_In(A_shift_out), .Load(Ld_B), .D(Bin),.A(Bout));
			
endmodule
